--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : MouseProject_modif                                           ==
--== Component : logisimTopLevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY logisimTopLevelShell IS
   PORT ( CLK_0      : IN  std_logic;
          PS_CLK_0   : IN  std_logic;
          PS_DATA_0  : IN  std_logic;
          REVERSE_0  : IN  std_logic;
          RST_0      : IN  std_logic;
          IS_LEFT_0  : OUT std_logic;
          n_ANODS_0  : OUT std_logic;
          n_ANODS_1  : OUT std_logic;
          n_ANODS_2  : OUT std_logic;
          n_ANODS_3  : OUT std_logic;
          n_CATODS_0 : OUT std_logic;
          n_CATODS_1 : OUT std_logic;
          n_CATODS_2 : OUT std_logic;
          n_CATODS_3 : OUT std_logic;
          n_CATODS_4 : OUT std_logic;
          n_CATODS_5 : OUT std_logic;
          n_CATODS_6 : OUT std_logic );
END ENTITY logisimTopLevelShell;
